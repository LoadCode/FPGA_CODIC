module rom (input clk,
                input wire [8:0] addr,
                output reg [31:0] data);

  //-- Memoria
  reg [31:0] angle_table [0:360];

  //-- Proceso de acceso a la memoria. 
  //-- Se ha elegido flanco de bajada en este ejemplo, pero
  //-- funciona igual si es de subida
  always @(posedge clk) begin
    data <= angle_table[addr];
  end

//-- Inicializacion de la memoria.
  initial begin
	angle_table[0] = 32'b00000000000000000000000000000000;
	angle_table[1] = 32'b00000000101101100000101101100001;
	angle_table[2] = 32'b00000001011011000001011011000001;
	angle_table[3] = 32'b00000010001000100010001000100010;
	angle_table[4] = 32'b00000010110110000010110110000011;
	angle_table[5] = 32'b00000011100011100011100011100100;
	angle_table[6] = 32'b00000100010001000100010001000100;
	angle_table[7] = 32'b00000100111110100100111110100101;
	angle_table[8] = 32'b00000101101100000101101100000110;
	angle_table[9] = 32'b00000110011001100110011001100110;
	angle_table[10] = 32'b00000111000111000111000111000111;
	angle_table[11] = 32'b00000111110100100111110100101000;
	angle_table[12] = 32'b00001000100010001000100010001001;
	angle_table[13] = 32'b00001001001111101001001111101001;
	angle_table[14] = 32'b00001001111101001001111101001010;
	angle_table[15] = 32'b00001010101010101010101010101011;
	angle_table[16] = 32'b00001011011000001011011000001011;
	angle_table[17] = 32'b00001100000101101100000101101100;
	angle_table[18] = 32'b00001100110011001100110011001101;
	angle_table[19] = 32'b00001101100000101101100000101110;
	angle_table[20] = 32'b00001110001110001110001110001110;
	angle_table[21] = 32'b00001110111011101110111011101111;
	angle_table[22] = 32'b00001111101001001111101001010000;
	angle_table[23] = 32'b00010000010110110000010110110000;
	angle_table[24] = 32'b00010001000100010001000100010001;
	angle_table[25] = 32'b00010001110001110001110001110010;
	angle_table[26] = 32'b00010010011111010010011111010010;
	angle_table[27] = 32'b00010011001100110011001100110011;
	angle_table[28] = 32'b00010011111010010011111010010100;
	angle_table[29] = 32'b00010100100111110100100111110101;
	angle_table[30] = 32'b00010101010101010101010101010101;
	angle_table[31] = 32'b00010110000010110110000010110110;
	angle_table[32] = 32'b00010110110000010110110000010111;
	angle_table[33] = 32'b00010111011101110111011101110111;
	angle_table[34] = 32'b00011000001011011000001011011000;
	angle_table[35] = 32'b00011000111000111000111000111001;
	angle_table[36] = 32'b00011001100110011001100110011010;
	angle_table[37] = 32'b00011010010011111010010011111010;
	angle_table[38] = 32'b00011011000001011011000001011011;
	angle_table[39] = 32'b00011011101110111011101110111100;
	angle_table[40] = 32'b00011100011100011100011100011100;
	angle_table[41] = 32'b00011101001001111101001001111101;
	angle_table[42] = 32'b00011101110111011101110111011110;
	angle_table[43] = 32'b00011110100100111110100100111111;
	angle_table[44] = 32'b00011111010010011111010010011111;
	angle_table[45] = 32'b00100000000000000000000000000000;
	angle_table[46] = 32'b00100000101101100000101101100001;
	angle_table[47] = 32'b00100001011011000001011011000001;
	angle_table[48] = 32'b00100010001000100010001000100010;
	angle_table[49] = 32'b00100010110110000010110110000011;
	angle_table[50] = 32'b00100011100011100011100011100100;
	angle_table[51] = 32'b00100100010001000100010001000100;
	angle_table[52] = 32'b00100100111110100100111110100101;
	angle_table[53] = 32'b00100101101100000101101100000110;
	angle_table[54] = 32'b00100110011001100110011001100110;
	angle_table[55] = 32'b00100111000111000111000111000111;
	angle_table[56] = 32'b00100111110100100111110100101000;
	angle_table[57] = 32'b00101000100010001000100010001001;
	angle_table[58] = 32'b00101001001111101001001111101001;
	angle_table[59] = 32'b00101001111101001001111101001010;
	angle_table[60] = 32'b00101010101010101010101010101011;
	angle_table[61] = 32'b00101011011000001011011000001011;
	angle_table[62] = 32'b00101100000101101100000101101100;
	angle_table[63] = 32'b00101100110011001100110011001101;
	angle_table[64] = 32'b00101101100000101101100000101110;
	angle_table[65] = 32'b00101110001110001110001110001110;
	angle_table[66] = 32'b00101110111011101110111011101111;
	angle_table[67] = 32'b00101111101001001111101001010000;
	angle_table[68] = 32'b00110000010110110000010110110000;
	angle_table[69] = 32'b00110001000100010001000100010001;
	angle_table[70] = 32'b00110001110001110001110001110010;
	angle_table[71] = 32'b00110010011111010010011111010010;
	angle_table[72] = 32'b00110011001100110011001100110011;
	angle_table[73] = 32'b00110011111010010011111010010100;
	angle_table[74] = 32'b00110100100111110100100111110101;
	angle_table[75] = 32'b00110101010101010101010101010101;
	angle_table[76] = 32'b00110110000010110110000010110110;
	angle_table[77] = 32'b00110110110000010110110000010111;
	angle_table[78] = 32'b00110111011101110111011101110111;
	angle_table[79] = 32'b00111000001011011000001011011000;
	angle_table[80] = 32'b00111000111000111000111000111001;
	angle_table[81] = 32'b00111001100110011001100110011010;
	angle_table[82] = 32'b00111010010011111010010011111010;
	angle_table[83] = 32'b00111011000001011011000001011011;
	angle_table[84] = 32'b00111011101110111011101110111100;
	angle_table[85] = 32'b00111100011100011100011100011100;
	angle_table[86] = 32'b00111101001001111101001001111101;
	angle_table[87] = 32'b00111101110111011101110111011110;
	angle_table[88] = 32'b00111110100100111110100100111111;
	angle_table[89] = 32'b00111111010010011111010010011111;
	angle_table[90] = 32'b01000000000000000000000000000000;
	angle_table[91] = 32'b01000000101101100000101101100001;
	angle_table[92] = 32'b01000001011011000001011011000001;
	angle_table[93] = 32'b01000010001000100010001000100010;
	angle_table[94] = 32'b01000010110110000010110110000011;
	angle_table[95] = 32'b01000011100011100011100011100100;
	angle_table[96] = 32'b01000100010001000100010001000100;
	angle_table[97] = 32'b01000100111110100100111110100101;
	angle_table[98] = 32'b01000101101100000101101100000110;
	angle_table[99] = 32'b01000110011001100110011001100110;
	angle_table[100] = 32'b01000111000111000111000111000111;
	angle_table[101] = 32'b01000111110100100111110100101000;
	angle_table[102] = 32'b01001000100010001000100010001001;
	angle_table[103] = 32'b01001001001111101001001111101001;
	angle_table[104] = 32'b01001001111101001001111101001010;
	angle_table[105] = 32'b01001010101010101010101010101011;
	angle_table[106] = 32'b01001011011000001011011000001011;
	angle_table[107] = 32'b01001100000101101100000101101100;
	angle_table[108] = 32'b01001100110011001100110011001101;
	angle_table[109] = 32'b01001101100000101101100000101110;
	angle_table[110] = 32'b01001110001110001110001110001110;
	angle_table[111] = 32'b01001110111011101110111011101111;
	angle_table[112] = 32'b01001111101001001111101001010000;
	angle_table[113] = 32'b01010000010110110000010110110000;
	angle_table[114] = 32'b01010001000100010001000100010001;
	angle_table[115] = 32'b01010001110001110001110001110010;
	angle_table[116] = 32'b01010010011111010010011111010010;
	angle_table[117] = 32'b01010011001100110011001100110011;
	angle_table[118] = 32'b01010011111010010011111010010100;
	angle_table[119] = 32'b01010100100111110100100111110101;
	angle_table[120] = 32'b01010101010101010101010101010101;
	angle_table[121] = 32'b01010110000010110110000010110110;
	angle_table[122] = 32'b01010110110000010110110000010111;
	angle_table[123] = 32'b01010111011101110111011101110111;
	angle_table[124] = 32'b01011000001011011000001011011000;
	angle_table[125] = 32'b01011000111000111000111000111001;
	angle_table[126] = 32'b01011001100110011001100110011010;
	angle_table[127] = 32'b01011010010011111010010011111010;
	angle_table[128] = 32'b01011011000001011011000001011011;
	angle_table[129] = 32'b01011011101110111011101110111100;
	angle_table[130] = 32'b01011100011100011100011100011100;
	angle_table[131] = 32'b01011101001001111101001001111101;
	angle_table[132] = 32'b01011101110111011101110111011110;
	angle_table[133] = 32'b01011110100100111110100100111111;
	angle_table[134] = 32'b01011111010010011111010010011111;
	angle_table[135] = 32'b01100000000000000000000000000000;
	angle_table[136] = 32'b01100000101101100000101101100001;
	angle_table[137] = 32'b01100001011011000001011011000001;
	angle_table[138] = 32'b01100010001000100010001000100010;
	angle_table[139] = 32'b01100010110110000010110110000011;
	angle_table[140] = 32'b01100011100011100011100011100100;
	angle_table[141] = 32'b01100100010001000100010001000100;
	angle_table[142] = 32'b01100100111110100100111110100101;
	angle_table[143] = 32'b01100101101100000101101100000110;
	angle_table[144] = 32'b01100110011001100110011001100110;
	angle_table[145] = 32'b01100111000111000111000111000111;
	angle_table[146] = 32'b01100111110100100111110100101000;
	angle_table[147] = 32'b01101000100010001000100010001001;
	angle_table[148] = 32'b01101001001111101001001111101001;
	angle_table[149] = 32'b01101001111101001001111101001010;
	angle_table[150] = 32'b01101010101010101010101010101011;
	angle_table[151] = 32'b01101011011000001011011000001011;
	angle_table[152] = 32'b01101100000101101100000101101100;
	angle_table[153] = 32'b01101100110011001100110011001101;
	angle_table[154] = 32'b01101101100000101101100000101110;
	angle_table[155] = 32'b01101110001110001110001110001110;
	angle_table[156] = 32'b01101110111011101110111011101111;
	angle_table[157] = 32'b01101111101001001111101001010000;
	angle_table[158] = 32'b01110000010110110000010110110000;
	angle_table[159] = 32'b01110001000100010001000100010001;
	angle_table[160] = 32'b01110001110001110001110001110010;
	angle_table[161] = 32'b01110010011111010010011111010010;
	angle_table[162] = 32'b01110011001100110011001100110011;
	angle_table[163] = 32'b01110011111010010011111010010100;
	angle_table[164] = 32'b01110100100111110100100111110101;
	angle_table[165] = 32'b01110101010101010101010101010101;
	angle_table[166] = 32'b01110110000010110110000010110110;
	angle_table[167] = 32'b01110110110000010110110000010111;
	angle_table[168] = 32'b01110111011101110111011101110111;
	angle_table[169] = 32'b01111000001011011000001011011000;
	angle_table[170] = 32'b01111000111000111000111000111001;
	angle_table[171] = 32'b01111001100110011001100110011010;
	angle_table[172] = 32'b01111010010011111010010011111010;
	angle_table[173] = 32'b01111011000001011011000001011011;
	angle_table[174] = 32'b01111011101110111011101110111100;
	angle_table[175] = 32'b01111100011100011100011100011100;
	angle_table[176] = 32'b01111101001001111101001001111101;
	angle_table[177] = 32'b01111101110111011101110111011110;
	angle_table[178] = 32'b01111110100100111110100100111111;
	angle_table[179] = 32'b01111111010010011111010010011111;
	angle_table[180] = 32'b10000000000000000000000000000000;
	angle_table[181] = 32'b10000000101101100000101101100001;
	angle_table[182] = 32'b10000001011011000001011011000001;
	angle_table[183] = 32'b10000010001000100010001000100010;
	angle_table[184] = 32'b10000010110110000010110110000011;
	angle_table[185] = 32'b10000011100011100011100011100100;
	angle_table[186] = 32'b10000100010001000100010001000100;
	angle_table[187] = 32'b10000100111110100100111110100101;
	angle_table[188] = 32'b10000101101100000101101100000110;
	angle_table[189] = 32'b10000110011001100110011001100110;
	angle_table[190] = 32'b10000111000111000111000111000111;
	angle_table[191] = 32'b10000111110100100111110100101000;
	angle_table[192] = 32'b10001000100010001000100010001001;
	angle_table[193] = 32'b10001001001111101001001111101001;
	angle_table[194] = 32'b10001001111101001001111101001010;
	angle_table[195] = 32'b10001010101010101010101010101011;
	angle_table[196] = 32'b10001011011000001011011000001011;
	angle_table[197] = 32'b10001100000101101100000101101100;
	angle_table[198] = 32'b10001100110011001100110011001101;
	angle_table[199] = 32'b10001101100000101101100000101110;
	angle_table[200] = 32'b10001110001110001110001110001110;
	angle_table[201] = 32'b10001110111011101110111011101111;
	angle_table[202] = 32'b10001111101001001111101001010000;
	angle_table[203] = 32'b10010000010110110000010110110000;
	angle_table[204] = 32'b10010001000100010001000100010001;
	angle_table[205] = 32'b10010001110001110001110001110010;
	angle_table[206] = 32'b10010010011111010010011111010010;
	angle_table[207] = 32'b10010011001100110011001100110011;
	angle_table[208] = 32'b10010011111010010011111010010100;
	angle_table[209] = 32'b10010100100111110100100111110101;
	angle_table[210] = 32'b10010101010101010101010101010101;
	angle_table[211] = 32'b10010110000010110110000010110110;
	angle_table[212] = 32'b10010110110000010110110000010111;
	angle_table[213] = 32'b10010111011101110111011101110111;
	angle_table[214] = 32'b10011000001011011000001011011000;
	angle_table[215] = 32'b10011000111000111000111000111001;
	angle_table[216] = 32'b10011001100110011001100110011010;
	angle_table[217] = 32'b10011010010011111010010011111010;
	angle_table[218] = 32'b10011011000001011011000001011011;
	angle_table[219] = 32'b10011011101110111011101110111100;
	angle_table[220] = 32'b10011100011100011100011100011100;
	angle_table[221] = 32'b10011101001001111101001001111101;
	angle_table[222] = 32'b10011101110111011101110111011110;
	angle_table[223] = 32'b10011110100100111110100100111111;
	angle_table[224] = 32'b10011111010010011111010010011111;
	angle_table[225] = 32'b10100000000000000000000000000000;
	angle_table[226] = 32'b10100000101101100000101101100001;
	angle_table[227] = 32'b10100001011011000001011011000001;
	angle_table[228] = 32'b10100010001000100010001000100010;
	angle_table[229] = 32'b10100010110110000010110110000011;
	angle_table[230] = 32'b10100011100011100011100011100100;
	angle_table[231] = 32'b10100100010001000100010001000100;
	angle_table[232] = 32'b10100100111110100100111110100101;
	angle_table[233] = 32'b10100101101100000101101100000110;
	angle_table[234] = 32'b10100110011001100110011001100110;
	angle_table[235] = 32'b10100111000111000111000111000111;
	angle_table[236] = 32'b10100111110100100111110100101000;
	angle_table[237] = 32'b10101000100010001000100010001001;
	angle_table[238] = 32'b10101001001111101001001111101001;
	angle_table[239] = 32'b10101001111101001001111101001010;
	angle_table[240] = 32'b10101010101010101010101010101011;
	angle_table[241] = 32'b10101011011000001011011000001011;
	angle_table[242] = 32'b10101100000101101100000101101100;
	angle_table[243] = 32'b10101100110011001100110011001101;
	angle_table[244] = 32'b10101101100000101101100000101110;
	angle_table[245] = 32'b10101110001110001110001110001110;
	angle_table[246] = 32'b10101110111011101110111011101111;
	angle_table[247] = 32'b10101111101001001111101001010000;
	angle_table[248] = 32'b10110000010110110000010110110000;
	angle_table[249] = 32'b10110001000100010001000100010001;
	angle_table[250] = 32'b10110001110001110001110001110010;
	angle_table[251] = 32'b10110010011111010010011111010010;
	angle_table[252] = 32'b10110011001100110011001100110011;
	angle_table[253] = 32'b10110011111010010011111010010100;
	angle_table[254] = 32'b10110100100111110100100111110101;
	angle_table[255] = 32'b10110101010101010101010101010101;
	angle_table[256] = 32'b10110110000010110110000010110110;
	angle_table[257] = 32'b10110110110000010110110000010111;
	angle_table[258] = 32'b10110111011101110111011101110111;
	angle_table[259] = 32'b10111000001011011000001011011000;
	angle_table[260] = 32'b10111000111000111000111000111001;
	angle_table[261] = 32'b10111001100110011001100110011010;
	angle_table[262] = 32'b10111010010011111010010011111010;
	angle_table[263] = 32'b10111011000001011011000001011011;
	angle_table[264] = 32'b10111011101110111011101110111100;
	angle_table[265] = 32'b10111100011100011100011100011100;
	angle_table[266] = 32'b10111101001001111101001001111101;
	angle_table[267] = 32'b10111101110111011101110111011110;
	angle_table[268] = 32'b10111110100100111110100100111111;
	angle_table[269] = 32'b10111111010010011111010010011111;
	angle_table[270] = 32'b11000000000000000000000000000000;
	angle_table[271] = 32'b11000000101101100000101101100001;
	angle_table[272] = 32'b11000001011011000001011011000001;
	angle_table[273] = 32'b11000010001000100010001000100010;
	angle_table[274] = 32'b11000010110110000010110110000011;
	angle_table[275] = 32'b11000011100011100011100011100100;
	angle_table[276] = 32'b11000100010001000100010001000100;
	angle_table[277] = 32'b11000100111110100100111110100101;
	angle_table[278] = 32'b11000101101100000101101100000110;
	angle_table[279] = 32'b11000110011001100110011001100110;
	angle_table[280] = 32'b11000111000111000111000111000111;
	angle_table[281] = 32'b11000111110100100111110100101000;
	angle_table[282] = 32'b11001000100010001000100010001001;
	angle_table[283] = 32'b11001001001111101001001111101001;
	angle_table[284] = 32'b11001001111101001001111101001010;
	angle_table[285] = 32'b11001010101010101010101010101011;
	angle_table[286] = 32'b11001011011000001011011000001011;
	angle_table[287] = 32'b11001100000101101100000101101100;
	angle_table[288] = 32'b11001100110011001100110011001101;
	angle_table[289] = 32'b11001101100000101101100000101110;
	angle_table[290] = 32'b11001110001110001110001110001110;
	angle_table[291] = 32'b11001110111011101110111011101111;
	angle_table[292] = 32'b11001111101001001111101001010000;
	angle_table[293] = 32'b11010000010110110000010110110000;
	angle_table[294] = 32'b11010001000100010001000100010001;
	angle_table[295] = 32'b11010001110001110001110001110010;
	angle_table[296] = 32'b11010010011111010010011111010010;
	angle_table[297] = 32'b11010011001100110011001100110011;
	angle_table[298] = 32'b11010011111010010011111010010100;
	angle_table[299] = 32'b11010100100111110100100111110101;
	angle_table[300] = 32'b11010101010101010101010101010101;
	angle_table[301] = 32'b11010110000010110110000010110110;
	angle_table[302] = 32'b11010110110000010110110000010111;
	angle_table[303] = 32'b11010111011101110111011101110111;
	angle_table[304] = 32'b11011000001011011000001011011000;
	angle_table[305] = 32'b11011000111000111000111000111001;
	angle_table[306] = 32'b11011001100110011001100110011010;
	angle_table[307] = 32'b11011010010011111010010011111010;
	angle_table[308] = 32'b11011011000001011011000001011011;
	angle_table[309] = 32'b11011011101110111011101110111100;
	angle_table[310] = 32'b11011100011100011100011100011100;
	angle_table[311] = 32'b11011101001001111101001001111101;
	angle_table[312] = 32'b11011101110111011101110111011110;
	angle_table[313] = 32'b11011110100100111110100100111111;
	angle_table[314] = 32'b11011111010010011111010010011111;
	angle_table[315] = 32'b11100000000000000000000000000000;
	angle_table[316] = 32'b11100000101101100000101101100001;
	angle_table[317] = 32'b11100001011011000001011011000001;
	angle_table[318] = 32'b11100010001000100010001000100010;
	angle_table[319] = 32'b11100010110110000010110110000011;
	angle_table[320] = 32'b11100011100011100011100011100100;
	angle_table[321] = 32'b11100100010001000100010001000100;
	angle_table[322] = 32'b11100100111110100100111110100101;
	angle_table[323] = 32'b11100101101100000101101100000110;
	angle_table[324] = 32'b11100110011001100110011001100110;
	angle_table[325] = 32'b11100111000111000111000111000111;
	angle_table[326] = 32'b11100111110100100111110100101000;
	angle_table[327] = 32'b11101000100010001000100010001001;
	angle_table[328] = 32'b11101001001111101001001111101001;
	angle_table[329] = 32'b11101001111101001001111101001010;
	angle_table[330] = 32'b11101010101010101010101010101011;
	angle_table[331] = 32'b11101011011000001011011000001011;
	angle_table[332] = 32'b11101100000101101100000101101100;
	angle_table[333] = 32'b11101100110011001100110011001101;
	angle_table[334] = 32'b11101101100000101101100000101110;
	angle_table[335] = 32'b11101110001110001110001110001110;
	angle_table[336] = 32'b11101110111011101110111011101111;
	angle_table[337] = 32'b11101111101001001111101001010000;
	angle_table[338] = 32'b11110000010110110000010110110000;
	angle_table[339] = 32'b11110001000100010001000100010001;
	angle_table[340] = 32'b11110001110001110001110001110010;
	angle_table[341] = 32'b11110010011111010010011111010010;
	angle_table[342] = 32'b11110011001100110011001100110011;
	angle_table[343] = 32'b11110011111010010011111010010100;
	angle_table[344] = 32'b11110100100111110100100111110101;
	angle_table[345] = 32'b11110101010101010101010101010101;
	angle_table[346] = 32'b11110110000010110110000010110110;
	angle_table[347] = 32'b11110110110000010110110000010111;
	angle_table[348] = 32'b11110111011101110111011101110111;
	angle_table[349] = 32'b11111000001011011000001011011000;
	angle_table[350] = 32'b11111000111000111000111000111001;
	angle_table[351] = 32'b11111001100110011001100110011010;
	angle_table[352] = 32'b11111010010011111010010011111010;
	angle_table[353] = 32'b11111011000001011011000001011011;
	angle_table[354] = 32'b11111011101110111011101110111100;
	angle_table[355] = 32'b11111100011100011100011100011100;
	angle_table[356] = 32'b11111101001001111101001001111101;
	angle_table[357] = 32'b11111101110111011101110111011110;
	angle_table[358] = 32'b11111110100100111110100100111111;
	angle_table[359] = 32'b11111111010010011111010010011111;
	
   end
	
endmodule
